// ----------------
// Project:
// ESA Elevator
// ----------------
//
// ----------------
// Group: 0
// 1234567: Wigald Boning
// 1234567: Oliver Dittrich 
// ----------------
//
// Description:
// ----------------
// elevator sensor interface
//

`timescale 1ns / 1ns

module sqrt

          (input wire         CLK,
           input wire         RESET,

           input wire         NEXT,
           input wire         PREVIOUS,

	   output reg 	      DONE,
	   output reg  [31:0] SQRT);
  
/* =============================INSERT CODE HERE======================================*/ 






/* ====================================================================================*/

endmodule 
